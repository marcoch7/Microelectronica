module map9v3 ( gnd, vdd, clock, reset, start, N, dp, done, counter, sr);

input gnd, vdd;
input clock;
input reset;
input start;
output done;
input [8:0] N;
output [8:0] dp;
output [7:0] counter;
output [7:0] sr;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_98__bF_buf3) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_98__bF_buf2) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_98__bF_buf1) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(_98_), .Y(_98__bF_buf0) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf4) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf3) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf2) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf1) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(clock), .Y(clock_bF_buf0) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_56__bF_buf4) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_56__bF_buf3) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_56__bF_buf2) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_56__bF_buf1) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(_56_), .Y(_56__bF_buf0) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(_97_), .Y(_97__bF_buf3) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(_97_), .Y(_97__bF_buf2) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_97_), .Y(_97__bF_buf1) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_97_), .Y(_97__bF_buf0) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .Y(_97_) );
	INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .Y(_98_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_117__3_), .B(_117__2_), .Y(_99_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_117__5_), .B(_117__4_), .Y(_100_) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_101_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_117__7_), .B(_117__6_), .Y(_102_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_117__1_), .B(_117__0_), .Y(_103_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_102_), .B(_103_), .Y(_104_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_101_), .Y(_105_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf3), .B(_105_), .C(_97__bF_buf3), .Y(_6_) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .Y(_106_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(state_1_), .Y(_107_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(startbuf_0_), .Y(_108_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(startbuf_1_), .B(_108_), .Y(_109_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_107_), .B(_109_), .C(_106_), .Y(_7_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_119__1_), .Y(_110_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .B(_97__bF_buf2), .C(_98__bF_buf2), .Y(_111_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_120__0_), .B(_111_), .Y(_112_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_110_), .B(_111_), .C(_112_), .Y(_2__1_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_119__2_), .Y(_113_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_120__1_), .Y(_114_) );
	MUX2X1 MUX2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_114_), .S(_111_), .Y(_2__2_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_119__3_), .Y(_115_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_120__2_), .Y(_116_) );
	MUX2X1 MUX2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .S(_111_), .Y(_2__3_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_119__4_), .Y(_8_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_120__3_), .Y(_9_) );
	MUX2X1 MUX2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_8_), .B(_9_), .S(_111_), .Y(_2__4_) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(_119__5_), .Y(_10_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(_120__4_), .Y(_11_) );
	MUX2X1 MUX2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_10_), .B(_11_), .S(_111_), .Y(_2__5_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(_119__6_), .Y(_12_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_120__5_), .Y(_13_) );
	MUX2X1 MUX2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_12_), .B(_13_), .S(_111_), .Y(_2__6_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_119__7_), .Y(_14_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_120__6_), .Y(_15_) );
	MUX2X1 MUX2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_14_), .B(_15_), .S(_111_), .Y(_2__7_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_119__8_), .Y(_16_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_120__7_), .Y(_17_) );
	MUX2X1 MUX2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_16_), .B(_17_), .S(_111_), .Y(_2__8_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_119__0_), .Y(_18_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(N[0]), .B(_111_), .Y(_19_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_18_), .B(_111_), .C(_19_), .Y(_2__0_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_120__5_), .B(_120__7_), .Y(_20_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_120__4_), .B(_9_), .Y(_21_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_120__3_), .B(_11_), .Y(_22_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_21_), .B(_22_), .C(_20_), .Y(_23_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_120__7_), .B(_13_), .Y(_24_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_120__5_), .B(_17_), .Y(_25_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_120__3_), .B(_120__4_), .Y(_26_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_24_), .B(_25_), .C(_26_), .Y(_27_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_23_), .B(_27_), .Y(_28_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_120__0_), .C(_97__bF_buf1), .Y(_29_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_28_), .B(state_3_), .C(_29_), .Y(_3__0_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_120__1_), .B(_98__bF_buf1), .C(_97__bF_buf0), .Y(_30_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf0), .B(_116_), .C(_30_), .Y(_3__2_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_120__2_), .B(_98__bF_buf3), .C(_97__bF_buf3), .Y(_31_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf2), .B(_9_), .C(_31_), .Y(_3__3_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_120__3_), .B(_98__bF_buf1), .C(_97__bF_buf2), .Y(_32_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf0), .B(_11_), .C(_32_), .Y(_3__4_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_120__4_), .B(_98__bF_buf3), .C(_97__bF_buf1), .Y(_33_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf2), .B(_13_), .C(_33_), .Y(_3__5_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_120__5_), .B(_98__bF_buf1), .C(_97__bF_buf0), .Y(_34_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf0), .B(_15_), .C(_34_), .Y(_3__6_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_120__6_), .B(_98__bF_buf3), .C(_97__bF_buf3), .Y(_35_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf2), .B(_17_), .C(_35_), .Y(_3__7_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(N[1]), .Y(_36_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(_117__0_), .B(_98__bF_buf1), .Y(_37_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf0), .B(_117__0_), .Y(_38_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_37_), .B(_38_), .C(_97__bF_buf2), .Y(_39_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_97__bF_buf1), .B(_36_), .C(_39_), .Y(_0__0_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(N[1]), .B(N[2]), .Y(_40_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(N[1]), .B(N[2]), .Y(_41_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_41_), .Y(_42_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_40_), .B(_42_), .C(state_0_), .Y(_43_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_103_), .B(state_3_), .Y(_44_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_117__1_), .Y(_45_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(_45_), .B(_37_), .Y(_46_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_44_), .B(_46_), .C(_97__bF_buf0), .Y(_47_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_43_), .B(_47_), .Y(_0__1_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_103_), .Y(_48_) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_117__2_), .Y(_49_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(N[3]), .Y(_50_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_41_), .Y(_51_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(N[3]), .B(_42_), .Y(_52_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_51_), .C(_52_), .Y(_53_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_49_), .C(_53_), .Y(_0__2_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(N[3]), .B(_42_), .C(N[4]), .Y(_54_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(N[4]), .Y(_55_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_50_), .B(_55_), .C(_41_), .Y(_57_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_54_), .Y(_58_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_117__3_), .B(_117__2_), .Y(_59_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_117__2_), .B(_48_), .C(_117__3_), .Y(_60_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_59_), .B(_48_), .C(_60_), .Y(_61_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_97__bF_buf3), .B(_61_), .Y(_62_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_97__bF_buf2), .B(_58_), .C(_62_), .Y(_0__3_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(N[5]), .Y(_63_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(N[3]), .B(N[4]), .Y(_64_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_64_), .B(_41_), .C(_63_), .Y(_65_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(N[5]), .B(_57_), .C(state_0_), .Y(_66_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_117__4_), .B(_59_), .Y(_67_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_44_), .Y(_68_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_44_), .C(_117__4_), .D(_68_), .Y(_69_) );
	OAI22X1 OAI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(_65_), .B(_66_), .C(state_0_), .D(_69_), .Y(_0__4_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(N[5]), .B(_57_), .C(N[6]), .Y(_70_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(N[5]), .B(N[6]), .Y(_71_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_57_), .B(_71_), .C(_70_), .Y(_72_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_101_), .Y(_73_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_117__5_), .Y(_74_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_67_), .B(_44_), .C(_74_), .Y(_75_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_75_), .C(_97__bF_buf1), .Y(_76_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_97__bF_buf0), .B(_72_), .C(_76_), .Y(_0__5_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(N[7]), .Y(_77_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(_71_), .B(_57_), .Y(_78_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_78_), .Y(_79_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(N[5]), .B(N[6]), .Y(_80_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_41_), .B(_64_), .C(_80_), .Y(_81_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(N[7]), .B(_81_), .C(state_0_), .Y(_82_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_117__6_), .Y(_83_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_99_), .B(_100_), .Y(_84_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(_83_), .B(_44_), .C(_84_), .Y(_85_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_48_), .B(_101_), .C(_117__6_), .Y(_86_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_85_), .B(_86_), .Y(_87_) );
	OAI22X1 OAI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_79_), .B(_82_), .C(state_0_), .D(_87_), .Y(_0__6_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(N[7]), .B(_81_), .C(N[8]), .Y(_88_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(N[8]), .Y(_89_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_77_), .B(_89_), .C(_78_), .Y(_90_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_88_), .C(_90_), .Y(_91_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(state_3_), .B(_105_), .C(_117__7_), .D(_85_), .Y(_92_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(state_0_), .B(_92_), .C(_91_), .Y(_0__7_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_118_), .Y(_93_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(state_2_), .Y(_94_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(state_4_), .B(_98__bF_buf3), .C(_94_), .Y(_95_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_93_), .C(state_0_), .Y(_1_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_120__0_), .B(_98__bF_buf2), .C(_97__bF_buf3), .Y(_96_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_98__bF_buf1), .B(_114_), .C(_96_), .Y(_3__1_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(state_1_), .Y(_4_) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_73_), .B(_102_), .Y(_5_) );
	INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(_56_) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_117__0_), .Y(counter[0]) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_117__1_), .Y(counter[1]) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_117__2_), .Y(counter[2]) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_117__3_), .Y(counter[3]) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_117__4_), .Y(counter[4]) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_117__5_), .Y(counter[5]) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_117__6_), .Y(counter[6]) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_117__7_), .Y(counter[7]) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_118_), .Y(done) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_119__0_), .Y(dp[0]) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_119__1_), .Y(dp[1]) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_119__2_), .Y(dp[2]) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_119__3_), .Y(dp[3]) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_119__4_), .Y(dp[4]) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_119__5_), .Y(dp[5]) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_119__6_), .Y(dp[6]) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_119__7_), .Y(dp[7]) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_119__8_), .Y(dp[8]) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_120__0_), .Y(sr[0]) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_120__1_), .Y(sr[1]) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_120__2_), .Y(sr[2]) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_120__3_), .Y(sr[3]) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_120__4_), .Y(sr[4]) );
	BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_120__5_), .Y(sr[5]) );
	BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_120__6_), .Y(sr[6]) );
	BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_120__7_), .Y(sr[7]) );
	DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_4_), .Q(state_0_), .R(vdd), .S(_56__bF_buf4) );
	DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_7_), .Q(state_1_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_5_), .Q(state_2_), .R(_56__bF_buf2), .S(vdd) );
	DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_6_), .Q(state_3_), .R(_56__bF_buf1), .S(vdd) );
	DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(state_2_), .Q(state_4_), .R(_56__bF_buf0), .S(vdd) );
	DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_2__0_), .Q(_119__0_), .R(_56__bF_buf4), .S(vdd) );
	DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_2__1_), .Q(_119__1_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_2__2_), .Q(_119__2_), .R(_56__bF_buf2), .S(vdd) );
	DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_2__3_), .Q(_119__3_), .R(_56__bF_buf1), .S(vdd) );
	DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_2__4_), .Q(_119__4_), .R(_56__bF_buf0), .S(vdd) );
	DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_2__5_), .Q(_119__5_), .R(_56__bF_buf4), .S(vdd) );
	DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_2__6_), .Q(_119__6_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_2__7_), .Q(_119__7_), .R(_56__bF_buf2), .S(vdd) );
	DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_2__8_), .Q(_119__8_), .R(_56__bF_buf1), .S(vdd) );
	DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_1_), .Q(_118_), .R(_56__bF_buf0), .S(vdd) );
	DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_0__0_), .Q(_117__0_), .R(_56__bF_buf4), .S(vdd) );
	DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_0__1_), .Q(_117__1_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_0__2_), .Q(_117__2_), .R(_56__bF_buf2), .S(vdd) );
	DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_0__3_), .Q(_117__3_), .R(_56__bF_buf1), .S(vdd) );
	DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_0__4_), .Q(_117__4_), .R(_56__bF_buf0), .S(vdd) );
	DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_0__5_), .Q(_117__5_), .R(_56__bF_buf4), .S(vdd) );
	DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_0__6_), .Q(_117__6_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_0__7_), .Q(_117__7_), .R(_56__bF_buf2), .S(vdd) );
	DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_3__0_), .Q(_120__0_), .R(_56__bF_buf1), .S(vdd) );
	DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_3__1_), .Q(_120__1_), .R(_56__bF_buf0), .S(vdd) );
	DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_3__2_), .Q(_120__2_), .R(_56__bF_buf4), .S(vdd) );
	DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(_3__3_), .Q(_120__3_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(_3__4_), .Q(_120__4_), .R(_56__bF_buf2), .S(vdd) );
	DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf1), .D(_3__5_), .Q(_120__5_), .R(_56__bF_buf1), .S(vdd) );
	DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf0), .D(_3__6_), .Q(_120__6_), .R(_56__bF_buf0), .S(vdd) );
	DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf4), .D(_3__7_), .Q(_120__7_), .R(_56__bF_buf4), .S(vdd) );
	DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf3), .D(start), .Q(startbuf_0_), .R(_56__bF_buf3), .S(vdd) );
	DFFSR DFFSR_33 ( .gnd(gnd), .vdd(vdd), .CLK(clock_bF_buf2), .D(startbuf_0_), .Q(startbuf_1_), .R(_56__bF_buf2), .S(vdd) );
endmodule
