module counter (clk, reset, enable, D, mode, Q, rco, load);

input clk;
input reset;
input enable;
output rco;
output load;
input [3:0] D;
input [1:0] mode;
output [3:0] Q;

wire vdd = 1'b1;
wire gnd = 1'b0;

	INVX1 INVX1_1 ( .A(reset), .Y(_2_) );
	INVX2 INVX2_1 ( .A(mode[1]), .Y(_3_) );
	INVX2 INVX2_2 ( .A(mode[0]), .Y(_4_) );
	NOR2X1 NOR2X1_1 ( .A(_3_), .B(_4_), .Y(_5_) );
	AND2X2 AND2X2_1 ( .A(_5_), .B(_2_), .Y(_1_) );
	NAND2X1 NAND2X1_1 ( .A(enable), .B(_2_), .Y(_6_) );
	NAND2X1 NAND2X1_2 ( .A(D[0]), .B(_5_), .Y(_7_) );
	INVX1 INVX1_2 ( .A(_36__0_), .Y(_8_) );
	OAI21X1 OAI21X1_1 ( .A(_3_), .B(_4_), .C(_8_), .Y(_9_) );
	AOI21X1 AOI21X1_1 ( .A(_7_), .B(_9_), .C(_6_), .Y(_0__0_) );
	NAND2X1 NAND2X1_3 ( .A(D[1]), .B(_5_), .Y(_10_) );
	XNOR2X1 XNOR2X1_1 ( .A(_36__0_), .B(_36__1_), .Y(_11_) );
	OAI21X1 OAI21X1_2 ( .A(mode[1]), .B(_4_), .C(_11_), .Y(_12_) );
	OAI21X1 OAI21X1_3 ( .A(_4_), .B(_11_), .C(_12_), .Y(_13_) );
	AOI21X1 AOI21X1_2 ( .A(_13_), .B(_10_), .C(_6_), .Y(_0__1_) );
	NOR2X1 NOR2X1_2 ( .A(mode[1]), .B(mode[0]), .Y(_14_) );
	AOI21X1 AOI21X1_3 ( .A(_36__0_), .B(_36__1_), .C(_36__2_), .Y(_15_) );
	INVX1 INVX1_3 ( .A(_15_), .Y(_16_) );
	NAND3X1 NAND3X1_1 ( .A(_36__0_), .B(_36__1_), .C(_36__2_), .Y(_17_) );
	AND2X2 AND2X2_2 ( .A(_16_), .B(_17_), .Y(_18_) );
	AOI22X1 AOI22X1_1 ( .A(D[2]), .B(_5_), .C(_14_), .D(_18_), .Y(_19_) );
	NOR2X1 NOR2X1_3 ( .A(mode[0]), .B(_3_), .Y(_20_) );
	NAND2X1 NAND2X1_4 ( .A(_17_), .B(_16_), .Y(_21_) );
	NAND2X1 NAND2X1_5 ( .A(mode[0]), .B(_3_), .Y(_22_) );
	INVX1 INVX1_4 ( .A(_36__2_), .Y(_23_) );
	NOR2X1 NOR2X1_4 ( .A(_36__0_), .B(_36__1_), .Y(_24_) );
	NAND2X1 NAND2X1_6 ( .A(_23_), .B(_24_), .Y(_25_) );
	OAI21X1 OAI21X1_4 ( .A(_36__0_), .B(_36__1_), .C(_36__2_), .Y(_26_) );
	AOI21X1 AOI21X1_4 ( .A(_25_), .B(_26_), .C(_22_), .Y(_27_) );
	AOI21X1 AOI21X1_5 ( .A(_20_), .B(_21_), .C(_27_), .Y(_28_) );
	AOI21X1 AOI21X1_6 ( .A(_19_), .B(_28_), .C(_6_), .Y(_0__2_) );
	XNOR2X1 XNOR2X1_2 ( .A(_17_), .B(_36__3_), .Y(_29_) );
	INVX1 INVX1_5 ( .A(_36__3_), .Y(_30_) );
	XNOR2X1 XNOR2X1_3 ( .A(_15_), .B(_30_), .Y(_31_) );
	AOI22X1 AOI22X1_2 ( .A(_29_), .B(_14_), .C(_20_), .D(_31_), .Y(_32_) );
	NAND3X1 NAND3X1_2 ( .A(_23_), .B(_36__3_), .C(_24_), .Y(_33_) );
	AOI21X1 AOI21X1_7 ( .A(_25_), .B(_30_), .C(_22_), .Y(_34_) );
	AOI22X1 AOI22X1_3 ( .A(D[3]), .B(_5_), .C(_33_), .D(_34_), .Y(_35_) );
	AOI21X1 AOI21X1_8 ( .A(_32_), .B(_35_), .C(_6_), .Y(_0__3_) );
	BUFX2 BUFX2_1 ( .A(_36__0_), .Y(Q[0]) );
	BUFX2 BUFX2_2 ( .A(_36__1_), .Y(Q[1]) );
	BUFX2 BUFX2_3 ( .A(_36__2_), .Y(Q[2]) );
	BUFX2 BUFX2_4 ( .A(_36__3_), .Y(Q[3]) );
	BUFX2 BUFX2_5 ( .A(_37_), .Y(load) );
	BUFX2 BUFX2_6 ( .A(gnd), .Y(rco) );
	DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_0__0_), .Q(_36__0_) );
	DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_0__1_), .Q(_36__1_) );
	DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_0__2_), .Q(_36__2_) );
	DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_0__3_), .Q(_36__3_) );
	DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_1_), .Q(_37_) );
endmodule
